library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;

entity ram is
port(clk, wr1, wr2 : in std_logic;
i, n : in std_logic_vector(3 downto 0);
j, set, sum : in std_logic_vector(7 downto 0);
y : out std_logic);
end ram;
architecture rtl of ram is
type ram_type is array (0 to 15, 0 to 255) of
std_logic;
type vec is array (0 to 255) of std_logic;
signal program: ram_type := (
    ('1', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0','0'),
    ('1', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0','0'),
    ('1', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0','0'),
    ('1', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0','0'),
    ('1', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0','0'),
    ('1', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0','0'),
    ('1', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0','0'),
    ('1', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0','0'),
    ('1', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0','0'),
    ('1', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0','0'),
    ('1', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0','0'),
    ('1', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0','0'),
    ('1', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0','0'),
    ('1', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0','0'),
    ('1', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0','0'),
    ('1', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0', '0','0', '0','0','0', '0','0','0', '0', '0','0','0','0', '0','0','0','0')
    
);
signal iminus1 : std_logic_vector(3 downto 0);
signal jminuss : std_logic_vector(7 downto 0);
signal s1, s2 : std_logic;

component sub is
    port (a, b : in std_logic_vector(7 downto 0);
    y : out std_logic_vector(7 downto 0));
end component;
component minus1 is
    port (a : in std_logic_vector(3 downto 0);
    y : out std_logic_vector(3 downto 0));
end component;

begin
s1 <= program(conv_integer(unsigned(iminus1)), conv_integer(unsigned(j)));
s2 <= program(conv_integer(unsigned(iminus1)), conv_integer(unsigned(jminuss)));
u1 : sub port map (j, set, jminuss);
u3 : minus1 port map (i, iminus1);
process(clk)
begin
if (rising_edge(clk)) then
if (wr1 = '1') then
program(conv_integer(unsigned(i)), conv_integer(unsigned(j))) <= s1;
elsif (wr2 = '1') then
program(conv_integer(unsigned(i)), conv_integer(unsigned(j))) <= s1 or s2;
end if;
end if;
end process;
y <= program(conv_integer(unsigned(n)), conv_integer(unsigned(sum)));
end rtl;